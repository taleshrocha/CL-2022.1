type byte is STD_LOGIC_VECTOR(0 to 7);
type barramento is ARRAY (0 down to 3) of byte;